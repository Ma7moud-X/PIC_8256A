library verilog;
use verilog.vl_types.all;
entity Data_bus_tb is
end Data_bus_tb;
