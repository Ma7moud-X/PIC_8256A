library verilog;
use verilog.vl_types.all;
entity Read_Write_Logic_tb is
end Read_Write_Logic_tb;
