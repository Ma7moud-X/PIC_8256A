library verilog;
use verilog.vl_types.all;
entity Control_Logic_tb is
end Control_Logic_tb;
