library verilog;
use verilog.vl_types.all;
entity IRR_tb is
end IRR_tb;
