library verilog;
use verilog.vl_types.all;
entity TOP_tb_1 is
end TOP_tb_1;
