library verilog;
use verilog.vl_types.all;
entity IMR_tb is
end IMR_tb;
