library verilog;
use verilog.vl_types.all;
entity ISR_tb is
end ISR_tb;
