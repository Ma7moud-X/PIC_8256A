library verilog;
use verilog.vl_types.all;
entity TOP_tb_2 is
end TOP_tb_2;
