library verilog;
use verilog.vl_types.all;
entity Priority_Resolver_tb is
end Priority_Resolver_tb;
