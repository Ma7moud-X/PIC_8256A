library verilog;
use verilog.vl_types.all;
entity Cascade_Buffer_tb is
end Cascade_Buffer_tb;
